library verilog;
use verilog.vl_types.all;
entity Common_Bus_System_vlg_vec_tst is
end Common_Bus_System_vlg_vec_tst;
