library verilog;
use verilog.vl_types.all;
entity ArithmaticLogicUnit_vlg_vec_tst is
end ArithmaticLogicUnit_vlg_vec_tst;
