library verilog;
use verilog.vl_types.all;
entity ShiftFunction_vlg_vec_tst is
end ShiftFunction_vlg_vec_tst;
